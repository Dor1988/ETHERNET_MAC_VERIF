typedef uvm_sequencer#(wb_tx) wb_proc_sqr;
