`include "eth_clockgen.v"
`include "eth_cop.v"
`include "eth_crc.v"
`include "eth_fifo.v"
`include "eth_maccontrol.v"
`include "ethmac_defines.v"
`include "eth_mac_rtl.svh"
`include "eth_macstatus.v"
`include "ethmac.v"
`include "eth_miim.v"
`include "eth_outputcontrol.v"
`include "eth_random.v"
`include "eth_receivecontrol.v"
`include "eth_registers.v"
`include "eth_register.v"
`include "eth_rxaddrcheck.v"
`include "eth_rxcounters.v"
`include "eth_rxethmac.v"
`include "eth_rxstatem.v"
`include "eth_shiftreg.v"
`include "eth_spram_256x32.v"
